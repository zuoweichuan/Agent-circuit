module mul12s_2PP ( A, B, O );
  input [11:0] A;
  input [11:0] B;
  output [23:0] O;

  wire [1344:0] N;

  assign N[0] = A[0] & B[0];
  assign N[1] = N[0];
  assign N[2] = A[0] & B[1];
  assign N[3] = N[2];
  assign N[4] = A[0] & B[2];
  assign N[5] = N[4];
  assign N[6] = A[0] & B[3];
  assign N[7] = N[6];
  assign N[8] = A[0] & B[4];
  assign N[9] = N[8];
  assign N[10] = A[0] & B[5];
  assign N[11] = N[10];
  assign N[12] = A[0] & B[6];
  assign N[13] = N[12];
  assign N[14] = A[0] & B[7];
  assign N[15] = N[14];
  assign N[16] = A[0] & B[8];
  assign N[17] = N[16];
  assign N[18] = A[0] & B[9];
  assign N[19] = N[18];
  assign N[20] = A[0] & B[10];
  assign N[21] = N[20];
  assign N[22] = A[0] & B[11];
  assign N[23] = ~N[22];
  assign N[24] = A[1] & B[0];
  assign N[25] = N[3] ^ N[24];
  assign N[26] = A[1] & B[0];
  assign N[27] = N[3] & N[26];
  assign N[28] = A[1] & B[1];
  assign N[29] = N[5] ^ N[28];
  assign N[30] = A[1] & B[1];
  assign N[31] = N[5] & N[30];
  assign N[32] = A[1] & B[2];
  assign N[33] = N[7] ^ N[32];
  assign N[34] = A[1] & B[2];
  assign N[35] = N[7] & N[34];
  assign N[36] = A[1] & B[3];
  assign N[37] = N[9] ^ N[36];
  assign N[38] = A[1] & B[3];
  assign N[39] = N[9] & N[38];
  assign N[40] = A[1] & B[4];
  assign N[41] = N[11] ^ N[40];
  assign N[42] = A[1] & B[4];
  assign N[43] = N[11] & N[42];
  assign N[44] = A[1] & B[5];
  assign N[45] = N[13] ^ N[44];
  assign N[46] = A[1] & B[5];
  assign N[47] = N[13] & N[46];
  assign N[48] = A[1] & B[6];
  assign N[49] = N[15] ^ N[48];
  assign N[50] = A[1] & B[6];
  assign N[51] = N[15] & N[50];
  assign N[52] = A[1] & B[7];
  assign N[53] = N[17] ^ N[52];
  assign N[54] = A[1] & B[7];
  assign N[55] = N[17] & N[54];
  assign N[56] = A[1] & B[8];
  assign N[57] = N[19] ^ N[56];
  assign N[58] = A[1] & B[8];
  assign N[59] = N[19] & N[58];
  assign N[60] = A[1] & B[9];
  assign N[61] = N[21] ^ N[60];
  assign N[62] = A[1] & B[9];
  assign N[63] = N[21] & N[62];
  assign N[64] = A[1] & B[10];
  assign N[65] = N[23] ^ N[64];
  assign N[66] = A[1] & B[10];
  assign N[67] = N[23] & N[66];
  assign N[68] = A[1] & B[11];
  assign N[69] = ~N[68];
  assign N[70] = 1'b1 ^  N[69];
  assign N[71] = A[1] & B[11];
  assign N[72] = ~N[71];
  assign N[73] = 1'b1 &  N[72];
  assign N[74] = N[29] ^ N[27];
  assign N[75] = A[2] & B[0];
  assign N[76] = N[74] ^ N[75];
  assign N[77] = N[29] & N[27];
  assign N[78] = A[2] & B[0];
  assign N[79] = A[2] & B[0];
  assign N[80] = N[27] & N[78];
  assign N[81] = N[29] & N[78];
  assign N[82] =  N[77] | N[80];
  assign N[83] = N[82] | N[81];
  assign N[84] = N[33] ^ N[31];
  assign N[85] = A[2] & B[1];
  assign N[86] = N[84] ^ N[85];
  assign N[87] = N[33] & N[31];
  assign N[88] = A[2] & B[1];
  assign N[89] = A[2] & B[1];
  assign N[90] = N[31] & N[88];
  assign N[91] = N[33] & N[88];
  assign N[92] =  N[87] | N[90];
  assign N[93] = N[92] | N[91];
  assign N[94] = N[37] ^ N[35];
  assign N[95] = A[2] & B[2];
  assign N[96] = N[94] ^ N[95];
  assign N[97] = N[37] & N[35];
  assign N[98] = A[2] & B[2];
  assign N[99] = A[2] & B[2];
  assign N[100] = N[35] & N[98];
  assign N[101] = N[37] & N[98];
  assign N[102] =  N[97] | N[100];
  assign N[103] = N[102] | N[101];
  assign N[104] = N[41] ^ N[39];
  assign N[105] = A[2] & B[3];
  assign N[106] = N[104] ^ N[105];
  assign N[107] = N[41] & N[39];
  assign N[108] = A[2] & B[3];
  assign N[109] = A[2] & B[3];
  assign N[110] = N[39] & N[108];
  assign N[111] = N[41] & N[108];
  assign N[112] =  N[107] | N[110];
  assign N[113] = N[112] | N[111];
  assign N[114] = N[45] ^ N[43];
  assign N[115] = A[2] & B[4];
  assign N[116] = N[114] ^ N[115];
  assign N[117] = N[45] & N[43];
  assign N[118] = A[2] & B[4];
  assign N[119] = A[2] & B[4];
  assign N[120] = N[43] & N[118];
  assign N[121] = N[45] & N[118];
  assign N[122] =  N[117] | N[120];
  assign N[123] = N[122] | N[121];
  assign N[124] = N[49] ^ N[47];
  assign N[125] = A[2] & B[5];
  assign N[126] = N[124] ^ N[125];
  assign N[127] = N[49] & N[47];
  assign N[128] = A[2] & B[5];
  assign N[129] = A[2] & B[5];
  assign N[130] = N[47] & N[128];
  assign N[131] = N[49] & N[128];
  assign N[132] =  N[127] | N[130];
  assign N[133] = N[132] | N[131];
  assign N[134] = N[53] ^ N[51];
  assign N[135] = A[2] & B[6];
  assign N[136] = N[134] ^ N[135];
  assign N[137] = N[53] & N[51];
  assign N[138] = A[2] & B[6];
  assign N[139] = A[2] & B[6];
  assign N[140] = N[51] & N[138];
  assign N[141] = N[53] & N[138];
  assign N[142] =  N[137] | N[140];
  assign N[143] = N[142] | N[141];
  assign N[144] = N[57] ^ N[55];
  assign N[145] = A[2] & B[7];
  assign N[146] = N[144] ^ N[145];
  assign N[147] = N[57] & N[55];
  assign N[148] = A[2] & B[7];
  assign N[149] = A[2] & B[7];
  assign N[150] = N[55] & N[148];
  assign N[151] = N[57] & N[148];
  assign N[152] =  N[147] | N[150];
  assign N[153] = N[152] | N[151];
  assign N[154] = N[61] ^ N[59];
  assign N[155] = A[2] & B[8];
  assign N[156] = N[154] ^ N[155];
  assign N[157] = N[61] & N[59];
  assign N[158] = A[2] & B[8];
  assign N[159] = A[2] & B[8];
  assign N[160] = N[59] & N[158];
  assign N[161] = N[61] & N[158];
  assign N[162] =  N[157] | N[160];
  assign N[163] = N[162] | N[161];
  assign N[164] = N[65] ^ N[63];
  assign N[165] = A[2] & B[9];
  assign N[166] = N[164] ^ N[165];
  assign N[167] = N[65] & N[63];
  assign N[168] = A[2] & B[9];
  assign N[169] = A[2] & B[9];
  assign N[170] = N[63] & N[168];
  assign N[171] = N[65] & N[168];
  assign N[172] =  N[167] | N[170];
  assign N[173] = N[172] | N[171];
  assign N[174] = N[70] ^ N[67];
  assign N[175] = A[2] & B[10];
  assign N[176] = N[174] ^ N[175];
  assign N[177] = N[70] & N[67];
  assign N[178] = A[2] & B[10];
  assign N[179] = A[2] & B[10];
  assign N[180] = N[67] & N[178];
  assign N[181] = N[70] & N[178];
  assign N[182] =  N[177] | N[180];
  assign N[183] = N[182] | N[181];
  assign N[184] = A[2] & B[11];
  assign N[185] = ~N[184];
  assign N[186] = N[73] ^  N[185];
  assign N[187] = A[2] & B[11];
  assign N[188] = ~N[187];
  assign N[189] = N[73] &  N[188];
  assign N[190] = N[86] ^ N[83];
  assign N[191] = A[3] & B[0];
  assign N[192] = N[190] ^ N[191];
  assign N[193] = N[86] & N[83];
  assign N[194] = A[3] & B[0];
  assign N[195] = A[3] & B[0];
  assign N[196] = N[83] & N[194];
  assign N[197] = N[86] & N[194];
  assign N[198] =  N[193] | N[196];
  assign N[199] = N[198] | N[197];
  assign N[200] = N[96] ^ N[93];
  assign N[201] = A[3] & B[1];
  assign N[202] = N[200] ^ N[201];
  assign N[203] = N[96] & N[93];
  assign N[204] = A[3] & B[1];
  assign N[205] = A[3] & B[1];
  assign N[206] = N[93] & N[204];
  assign N[207] = N[96] & N[204];
  assign N[208] =  N[203] | N[206];
  assign N[209] = N[208] | N[207];
  assign N[210] = N[106] ^ N[103];
  assign N[211] = A[3] & B[2];
  assign N[212] = N[210] ^ N[211];
  assign N[213] = N[106] & N[103];
  assign N[214] = A[3] & B[2];
  assign N[215] = A[3] & B[2];
  assign N[216] = N[103] & N[214];
  assign N[217] = N[106] & N[214];
  assign N[218] =  N[213] | N[216];
  assign N[219] = N[218] | N[217];
  assign N[220] = N[116] ^ N[113];
  assign N[221] = A[3] & B[3];
  assign N[222] = N[220] ^ N[221];
  assign N[223] = N[116] & N[113];
  assign N[224] = A[3] & B[3];
  assign N[225] = A[3] & B[3];
  assign N[226] = N[113] & N[224];
  assign N[227] = N[116] & N[224];
  assign N[228] =  N[223] | N[226];
  assign N[229] = N[228] | N[227];
  assign N[230] = N[126] ^ N[123];
  assign N[231] = A[3] & B[4];
  assign N[232] = N[230] ^ N[231];
  assign N[233] = N[126] & N[123];
  assign N[234] = A[3] & B[4];
  assign N[235] = A[3] & B[4];
  assign N[236] = N[123] & N[234];
  assign N[237] = N[126] & N[234];
  assign N[238] =  N[233] | N[236];
  assign N[239] = N[238] | N[237];
  assign N[240] = N[136] ^ N[133];
  assign N[241] = A[3] & B[5];
  assign N[242] = N[240] ^ N[241];
  assign N[243] = N[136] & N[133];
  assign N[244] = A[3] & B[5];
  assign N[245] = A[3] & B[5];
  assign N[246] = N[133] & N[244];
  assign N[247] = N[136] & N[244];
  assign N[248] =  N[243] | N[246];
  assign N[249] = N[248] | N[247];
  assign N[250] = N[146] ^ N[143];
  assign N[251] = A[3] & B[6];
  assign N[252] = N[250] ^ N[251];
  assign N[253] = N[146] & N[143];
  assign N[254] = A[3] & B[6];
  assign N[255] = A[3] & B[6];
  assign N[256] = N[143] & N[254];
  assign N[257] = N[146] & N[254];
  assign N[258] =  N[253] | N[256];
  assign N[259] = N[258] | N[257];
  assign N[260] = N[156] ^ N[153];
  assign N[261] = A[3] & B[7];
  assign N[262] = N[260] ^ N[261];
  assign N[263] = N[156] & N[153];
  assign N[264] = A[3] & B[7];
  assign N[265] = A[3] & B[7];
  assign N[266] = N[153] & N[264];
  assign N[267] = N[156] & N[264];
  assign N[268] =  N[263] | N[266];
  assign N[269] = N[268] | N[267];
  assign N[270] = N[166] ^ N[163];
  assign N[271] = A[3] & B[8];
  assign N[272] = N[270] ^ N[271];
  assign N[273] = N[166] & N[163];
  assign N[274] = A[3] & B[8];
  assign N[275] = A[3] & B[8];
  assign N[276] = N[163] & N[274];
  assign N[277] = N[166] & N[274];
  assign N[278] =  N[273] | N[276];
  assign N[279] = N[278] | N[277];
  assign N[280] = N[176] ^ N[173];
  assign N[281] = A[3] & B[9];
  assign N[282] = N[280] ^ N[281];
  assign N[283] = N[176] & N[173];
  assign N[284] = A[3] & B[9];
  assign N[285] = A[3] & B[9];
  assign N[286] = N[173] & N[284];
  assign N[287] = N[176] & N[284];
  assign N[288] =  N[283] | N[286];
  assign N[289] = N[288] | N[287];
  assign N[290] = N[186] ^ N[183];
  assign N[291] = A[3] & B[10];
  assign N[292] = N[290] ^ N[291];
  assign N[293] = N[186] & N[183];
  assign N[294] = A[3] & B[10];
  assign N[295] = A[3] & B[10];
  assign N[296] = N[183] & N[294];
  assign N[297] = N[186] & N[294];
  assign N[298] =  N[293] | N[296];
  assign N[299] = N[298] | N[297];
  assign N[300] = A[3] & B[11];
  assign N[301] = ~N[300];
  assign N[302] = N[189] ^  N[301];
  assign N[303] = A[3] & B[11];
  assign N[304] = ~N[303];
  assign N[305] = N[189] &  N[304];
  assign N[306] = N[202] ^ N[199];
  assign N[307] = A[4] & B[0];
  assign N[308] = N[306] ^ N[307];
  assign N[309] = N[202] & N[199];
  assign N[310] = A[4] & B[0];
  assign N[311] = A[4] & B[0];
  assign N[312] = N[199] & N[310];
  assign N[313] = N[202] & N[310];
  assign N[314] =  N[309] | N[312];
  assign N[315] = N[314] | N[313];
  assign N[316] = N[212] ^ N[209];
  assign N[317] = A[4] & B[1];
  assign N[318] = N[316] ^ N[317];
  assign N[319] = N[212] & N[209];
  assign N[320] = A[4] & B[1];
  assign N[321] = A[4] & B[1];
  assign N[322] = N[209] & N[320];
  assign N[323] = N[212] & N[320];
  assign N[324] =  N[319] | N[322];
  assign N[325] = N[324] | N[323];
  assign N[326] = N[222] ^ N[219];
  assign N[327] = A[4] & B[2];
  assign N[328] = N[326] ^ N[327];
  assign N[329] = N[222] & N[219];
  assign N[330] = A[4] & B[2];
  assign N[331] = A[4] & B[2];
  assign N[332] = N[219] & N[330];
  assign N[333] = N[222] & N[330];
  assign N[334] =  N[329] | N[332];
  assign N[335] = N[334] | N[333];
  assign N[336] = N[232] ^ N[229];
  assign N[337] = A[4] & B[3];
  assign N[338] = N[336] ^ N[337];
  assign N[339] = N[232] & N[229];
  assign N[340] = A[4] & B[3];
  assign N[341] = A[4] & B[3];
  assign N[342] = N[229] & N[340];
  assign N[343] = N[232] & N[340];
  assign N[344] =  N[339] | N[342];
  assign N[345] = N[344] | N[343];
  assign N[346] = N[242] ^ N[239];
  assign N[347] = A[4] & B[4];
  assign N[348] = N[346] ^ N[347];
  assign N[349] = N[242] & N[239];
  assign N[350] = A[4] & B[4];
  assign N[351] = A[4] & B[4];
  assign N[352] = N[239] & N[350];
  assign N[353] = N[242] & N[350];
  assign N[354] =  N[349] | N[352];
  assign N[355] = N[354] | N[353];
  assign N[356] = N[252] ^ N[249];
  assign N[357] = A[4] & B[5];
  assign N[358] = N[356] ^ N[357];
  assign N[359] = N[252] & N[249];
  assign N[360] = A[4] & B[5];
  assign N[361] = A[4] & B[5];
  assign N[362] = N[249] & N[360];
  assign N[363] = N[252] & N[360];
  assign N[364] =  N[359] | N[362];
  assign N[365] = N[364] | N[363];
  assign N[366] = N[262] ^ N[259];
  assign N[367] = A[4] & B[6];
  assign N[368] = N[366] ^ N[367];
  assign N[369] = N[262] & N[259];
  assign N[370] = A[4] & B[6];
  assign N[371] = A[4] & B[6];
  assign N[372] = N[259] & N[370];
  assign N[373] = N[262] & N[370];
  assign N[374] =  N[369] | N[372];
  assign N[375] = N[374] | N[373];
  assign N[376] = N[272] ^ N[269];
  assign N[377] = A[4] & B[7];
  assign N[378] = N[376] ^ N[377];
  assign N[379] = N[272] & N[269];
  assign N[380] = A[4] & B[7];
  assign N[381] = A[4] & B[7];
  assign N[382] = N[269] & N[380];
  assign N[383] = N[272] & N[380];
  assign N[384] =  N[379] | N[382];
  assign N[385] = N[384] | N[383];
  assign N[386] = N[282] ^ N[279];
  assign N[387] = A[4] & B[8];
  assign N[388] = N[386] ^ N[387];
  assign N[389] = N[282] & N[279];
  assign N[390] = A[4] & B[8];
  assign N[391] = A[4] & B[8];
  assign N[392] = N[279] & N[390];
  assign N[393] = N[282] & N[390];
  assign N[394] =  N[389] | N[392];
  assign N[395] = N[394] | N[393];
  assign N[396] = N[292] ^ N[289];
  assign N[397] = A[4] & B[9];
  assign N[398] = N[396] ^ N[397];
  assign N[399] = N[292] & N[289];
  assign N[400] = A[4] & B[9];
  assign N[401] = A[4] & B[9];
  assign N[402] = N[289] & N[400];
  assign N[403] = N[292] & N[400];
  assign N[404] =  N[399] | N[402];
  assign N[405] = N[404] | N[403];
  assign N[406] = N[302] ^ N[299];
  assign N[407] = A[4] & B[10];
  assign N[408] = N[406] ^ N[407];
  assign N[409] = N[302] & N[299];
  assign N[410] = A[4] & B[10];
  assign N[411] = A[4] & B[10];
  assign N[412] = N[299] & N[410];
  assign N[413] = N[302] & N[410];
  assign N[414] =  N[409] | N[412];
  assign N[415] = N[414] | N[413];
  assign N[416] = A[4] & B[11];
  assign N[417] = ~N[416];
  assign N[418] = N[305] ^  N[417];
  assign N[419] = A[4] & B[11];
  assign N[420] = ~N[419];
  assign N[421] = N[305] &  N[420];
  assign N[422] = N[318] ^ N[315];
  assign N[423] = A[5] & B[0];
  assign N[424] = N[422] ^ N[423];
  assign N[425] = N[318] & N[315];
  assign N[426] = A[5] & B[0];
  assign N[427] = A[5] & B[0];
  assign N[428] = N[315] & N[426];
  assign N[429] = N[318] & N[426];
  assign N[430] =  N[425] | N[428];
  assign N[431] = N[430] | N[429];
  assign N[432] = N[328] ^ N[325];
  assign N[433] = A[5] & B[1];
  assign N[434] = N[432] ^ N[433];
  assign N[435] = N[328] & N[325];
  assign N[436] = A[5] & B[1];
  assign N[437] = A[5] & B[1];
  assign N[438] = N[325] & N[436];
  assign N[439] = N[328] & N[436];
  assign N[440] =  N[435] | N[438];
  assign N[441] = N[440] | N[439];
  assign N[442] = N[338] ^ N[335];
  assign N[443] = A[5] & B[2];
  assign N[444] = N[442] ^ N[443];
  assign N[445] = N[338] & N[335];
  assign N[446] = A[5] & B[2];
  assign N[447] = A[5] & B[2];
  assign N[448] = N[335] & N[446];
  assign N[449] = N[338] & N[446];
  assign N[450] =  N[445] | N[448];
  assign N[451] = N[450] | N[449];
  assign N[452] = N[348] ^ N[345];
  assign N[453] = A[5] & B[3];
  assign N[454] = N[452] ^ N[453];
  assign N[455] = N[348] & N[345];
  assign N[456] = A[5] & B[3];
  assign N[457] = A[5] & B[3];
  assign N[458] = N[345] & N[456];
  assign N[459] = N[348] & N[456];
  assign N[460] =  N[455] | N[458];
  assign N[461] = N[460] | N[459];
  assign N[462] = N[358] ^ N[355];
  assign N[463] = A[5] & B[4];
  assign N[464] = N[462] ^ N[463];
  assign N[465] = N[358] & N[355];
  assign N[466] = A[5] & B[4];
  assign N[467] = A[5] & B[4];
  assign N[468] = N[355] & N[466];
  assign N[469] = N[358] & N[466];
  assign N[470] =  N[465] | N[468];
  assign N[471] = N[470] | N[469];
  assign N[472] = N[368] ^ N[365];
  assign N[473] = A[5] & B[5];
  assign N[474] = N[472] ^ N[473];
  assign N[475] = N[368] & N[365];
  assign N[476] = A[5] & B[5];
  assign N[477] = A[5] & B[5];
  assign N[478] = N[365] & N[476];
  assign N[479] = N[368] & N[476];
  assign N[480] =  N[475] | N[478];
  assign N[481] = N[480] | N[479];
  assign N[482] = N[378] ^ N[375];
  assign N[483] = A[5] & B[6];
  assign N[484] = N[482] ^ N[483];
  assign N[485] = N[378] & N[375];
  assign N[486] = A[5] & B[6];
  assign N[487] = A[5] & B[6];
  assign N[488] = N[375] & N[486];
  assign N[489] = N[378] & N[486];
  assign N[490] =  N[485] | N[488];
  assign N[491] = N[490] | N[489];
  assign N[492] = N[388] ^ N[385];
  assign N[493] = A[5] & B[7];
  assign N[494] = N[492] ^ N[493];
  assign N[495] = N[388] & N[385];
  assign N[496] = A[5] & B[7];
  assign N[497] = A[5] & B[7];
  assign N[498] = N[385] & N[496];
  assign N[499] = N[388] & N[496];
  assign N[500] =  N[495] | N[498];
  assign N[501] = N[500] | N[499];
  assign N[502] = N[398] ^ N[395];
  assign N[503] = A[5] & B[8];
  assign N[504] = N[502] ^ N[503];
  assign N[505] = N[398] & N[395];
  assign N[506] = A[5] & B[8];
  assign N[507] = A[5] & B[8];
  assign N[508] = N[395] & N[506];
  assign N[509] = N[398] & N[506];
  assign N[510] =  N[505] | N[508];
  assign N[511] = N[510] | N[509];
  assign N[512] = N[408] ^ N[405];
  assign N[513] = A[5] & B[9];
  assign N[514] = N[512] ^ N[513];
  assign N[515] = N[408] & N[405];
  assign N[516] = A[5] & B[9];
  assign N[517] = A[5] & B[9];
  assign N[518] = N[405] & N[516];
  assign N[519] = N[408] & N[516];
  assign N[520] =  N[515] | N[518];
  assign N[521] = N[520] | N[519];
  assign N[522] = N[418] ^ N[415];
  assign N[523] = A[5] & B[10];
  assign N[524] = N[522] ^ N[523];
  assign N[525] = N[418] & N[415];
  assign N[526] = A[5] & B[10];
  assign N[527] = A[5] & B[10];
  assign N[528] = N[415] & N[526];
  assign N[529] = N[418] & N[526];
  assign N[530] =  N[525] | N[528];
  assign N[531] = N[530] | N[529];
  assign N[532] = A[5] & B[11];
  assign N[533] = ~N[532];
  assign N[534] = N[421] ^  N[533];
  assign N[535] = A[5] & B[11];
  assign N[536] = ~N[535];
  assign N[537] = N[421] &  N[536];
  assign N[538] = N[434] ^ N[431];
  assign N[539] = A[6] & B[0];
  assign N[540] = N[538] ^ N[539];
  assign N[541] = N[434] & N[431];
  assign N[542] = A[6] & B[0];
  assign N[543] = A[6] & B[0];
  assign N[544] = N[431] & N[542];
  assign N[545] = N[434] & N[542];
  assign N[546] =  N[541] | N[544];
  assign N[547] = N[546] | N[545];
  assign N[548] = N[444] ^ N[441];
  assign N[549] = A[6] & B[1];
  assign N[550] = N[548] ^ N[549];
  assign N[551] = N[444] & N[441];
  assign N[552] = A[6] & B[1];
  assign N[553] = A[6] & B[1];
  assign N[554] = N[441] & N[552];
  assign N[555] = N[444] & N[552];
  assign N[556] =  N[551] | N[554];
  assign N[557] = N[556] | N[555];
  assign N[558] = N[454] ^ N[451];
  assign N[559] = A[6] & B[2];
  assign N[560] = N[558] ^ N[559];
  assign N[561] = N[454] & N[451];
  assign N[562] = A[6] & B[2];
  assign N[563] = A[6] & B[2];
  assign N[564] = N[451] & N[562];
  assign N[565] = N[454] & N[562];
  assign N[566] =  N[561] | N[564];
  assign N[567] = N[566] | N[565];
  assign N[568] = N[464] ^ N[461];
  assign N[569] = A[6] & B[3];
  assign N[570] = N[568] ^ N[569];
  assign N[571] = N[464] & N[461];
  assign N[572] = A[6] & B[3];
  assign N[573] = A[6] & B[3];
  assign N[574] = N[461] & N[572];
  assign N[575] = N[464] & N[572];
  assign N[576] =  N[571] | N[574];
  assign N[577] = N[576] | N[575];
  assign N[578] = N[474] ^ N[471];
  assign N[579] = A[6] & B[4];
  assign N[580] = N[578] ^ N[579];
  assign N[581] = N[474] & N[471];
  assign N[582] = A[6] & B[4];
  assign N[583] = A[6] & B[4];
  assign N[584] = N[471] & N[582];
  assign N[585] = N[474] & N[582];
  assign N[586] =  N[581] | N[584];
  assign N[587] = N[586] | N[585];
  assign N[588] = N[484] ^ N[481];
  assign N[589] = A[6] & B[5];
  assign N[590] = N[588] ^ N[589];
  assign N[591] = N[484] & N[481];
  assign N[592] = A[6] & B[5];
  assign N[593] = A[6] & B[5];
  assign N[594] = N[481] & N[592];
  assign N[595] = N[484] & N[592];
  assign N[596] =  N[591] | N[594];
  assign N[597] = N[596] | N[595];
  assign N[598] = N[494] ^ N[491];
  assign N[599] = A[6] & B[6];
  assign N[600] = N[598] ^ N[599];
  assign N[601] = N[494] & N[491];
  assign N[602] = A[6] & B[6];
  assign N[603] = A[6] & B[6];
  assign N[604] = N[491] & N[602];
  assign N[605] = N[494] & N[602];
  assign N[606] =  N[601] | N[604];
  assign N[607] = N[606] | N[605];
  assign N[608] = N[504] ^ N[501];
  assign N[609] = A[6] & B[7];
  assign N[610] = N[608] ^ N[609];
  assign N[611] = N[504] & N[501];
  assign N[612] = A[6] & B[7];
  assign N[613] = A[6] & B[7];
  assign N[614] = N[501] & N[612];
  assign N[615] = N[504] & N[612];
  assign N[616] =  N[611] | N[614];
  assign N[617] = N[616] | N[615];
  assign N[618] = N[514] ^ N[511];
  assign N[619] = A[6] & B[8];
  assign N[620] = N[618] ^ N[619];
  assign N[621] = N[514] & N[511];
  assign N[622] = A[6] & B[8];
  assign N[623] = A[6] & B[8];
  assign N[624] = N[511] & N[622];
  assign N[625] = N[514] & N[622];
  assign N[626] =  N[621] | N[624];
  assign N[627] = N[626] | N[625];
  assign N[628] = N[524] ^ N[521];
  assign N[629] = A[6] & B[9];
  assign N[630] = N[628] ^ N[629];
  assign N[631] = N[524] & N[521];
  assign N[632] = A[6] & B[9];
  assign N[633] = A[6] & B[9];
  assign N[634] = N[521] & N[632];
  assign N[635] = N[524] & N[632];
  assign N[636] =  N[631] | N[634];
  assign N[637] = N[636] | N[635];
  assign N[638] = N[534] ^ N[531];
  assign N[639] = A[6] & B[10];
  assign N[640] = N[638] ^ N[639];
  assign N[641] = N[534] & N[531];
  assign N[642] = A[6] & B[10];
  assign N[643] = A[6] & B[10];
  assign N[644] = N[531] & N[642];
  assign N[645] = N[534] & N[642];
  assign N[646] =  N[641] | N[644];
  assign N[647] = N[646] | N[645];
  assign N[648] = A[6] & B[11];
  assign N[649] = ~N[648];
  assign N[650] = N[537] ^  N[649];
  assign N[651] = A[6] & B[11];
  assign N[652] = ~N[651];
  assign N[653] = N[537] &  N[652];
  assign N[654] = N[550] ^ N[547];
  assign N[655] = A[7] & B[0];
  assign N[656] = N[654] ^ N[655];
  assign N[657] = N[550] & N[547];
  assign N[658] = A[7] & B[0];
  assign N[659] = A[7] & B[0];
  assign N[660] = N[547] & N[658];
  assign N[661] = N[550] & N[658];
  assign N[662] =  N[657] | N[660];
  assign N[663] = N[662] | N[661];
  assign N[664] = N[560] ^ N[557];
  assign N[665] = A[7] & B[1];
  assign N[666] = N[664] ^ N[665];
  assign N[667] = N[560] & N[557];
  assign N[668] = A[7] & B[1];
  assign N[669] = A[7] & B[1];
  assign N[670] = N[557] & N[668];
  assign N[671] = N[560] & N[668];
  assign N[672] =  N[667] | N[670];
  assign N[673] = N[672] | N[671];
  assign N[674] = N[570] ^ N[567];
  assign N[675] = A[7] & B[2];
  assign N[676] = N[674] ^ N[675];
  assign N[677] = N[570] & N[567];
  assign N[678] = A[7] & B[2];
  assign N[679] = A[7] & B[2];
  assign N[680] = N[567] & N[678];
  assign N[681] = N[570] & N[678];
  assign N[682] =  N[677] | N[680];
  assign N[683] = N[682] | N[681];
  assign N[684] = N[580] ^ N[577];
  assign N[685] = A[7] & B[3];
  assign N[686] = N[684] ^ N[685];
  assign N[687] = N[580] & N[577];
  assign N[688] = A[7] & B[3];
  assign N[689] = A[7] & B[3];
  assign N[690] = N[577] & N[688];
  assign N[691] = N[580] & N[688];
  assign N[692] =  N[687] | N[690];
  assign N[693] = N[692] | N[691];
  assign N[694] = N[590] ^ N[587];
  assign N[695] = A[7] & B[4];
  assign N[696] = N[694] ^ N[695];
  assign N[697] = N[590] & N[587];
  assign N[698] = A[7] & B[4];
  assign N[699] = A[7] & B[4];
  assign N[700] = N[587] & N[698];
  assign N[701] = N[590] & N[698];
  assign N[702] =  N[697] | N[700];
  assign N[703] = N[702] | N[701];
  assign N[704] = N[600] ^ N[597];
  assign N[705] = A[7] & B[5];
  assign N[706] = N[704] ^ N[705];
  assign N[707] = N[600] & N[597];
  assign N[708] = A[7] & B[5];
  assign N[709] = A[7] & B[5];
  assign N[710] = N[597] & N[708];
  assign N[711] = N[600] & N[708];
  assign N[712] =  N[707] | N[710];
  assign N[713] = N[712] | N[711];
  assign N[714] = N[610] ^ N[607];
  assign N[715] = A[7] & B[6];
  assign N[716] = N[714] ^ N[715];
  assign N[717] = N[610] & N[607];
  assign N[718] = A[7] & B[6];
  assign N[719] = A[7] & B[6];
  assign N[720] = N[607] & N[718];
  assign N[721] = N[610] & N[718];
  assign N[722] =  N[717] | N[720];
  assign N[723] = N[722] | N[721];
  assign N[724] = N[620] ^ N[617];
  assign N[725] = A[7] & B[7];
  assign N[726] = N[724] ^ N[725];
  assign N[727] = N[620] & N[617];
  assign N[728] = A[7] & B[7];
  assign N[729] = A[7] & B[7];
  assign N[730] = N[617] & N[728];
  assign N[731] = N[620] & N[728];
  assign N[732] =  N[727] | N[730];
  assign N[733] = N[732] | N[731];
  assign N[734] = N[630] ^ N[627];
  assign N[735] = A[7] & B[8];
  assign N[736] = N[734] ^ N[735];
  assign N[737] = N[630] & N[627];
  assign N[738] = A[7] & B[8];
  assign N[739] = A[7] & B[8];
  assign N[740] = N[627] & N[738];
  assign N[741] = N[630] & N[738];
  assign N[742] =  N[737] | N[740];
  assign N[743] = N[742] | N[741];
  assign N[744] = N[640] ^ N[637];
  assign N[745] = A[7] & B[9];
  assign N[746] = N[744] ^ N[745];
  assign N[747] = N[640] & N[637];
  assign N[748] = A[7] & B[9];
  assign N[749] = A[7] & B[9];
  assign N[750] = N[637] & N[748];
  assign N[751] = N[640] & N[748];
  assign N[752] =  N[747] | N[750];
  assign N[753] = N[752] | N[751];
  assign N[754] = N[650] ^ N[647];
  assign N[755] = A[7] & B[10];
  assign N[756] = N[754] ^ N[755];
  assign N[757] = N[650] & N[647];
  assign N[758] = A[7] & B[10];
  assign N[759] = A[7] & B[10];
  assign N[760] = N[647] & N[758];
  assign N[761] = N[650] & N[758];
  assign N[762] =  N[757] | N[760];
  assign N[763] = N[762] | N[761];
  assign N[764] = A[7] & B[11];
  assign N[765] = ~N[764];
  assign N[766] = N[653] ^  N[765];
  assign N[767] = A[7] & B[11];
  assign N[768] = ~N[767];
  assign N[769] = N[653] &  N[768];
  assign N[770] = N[666] ^ N[663];
  assign N[771] = A[8] & B[0];
  assign N[772] = N[770] ^ N[771];
  assign N[773] = N[666] & N[663];
  assign N[774] = A[8] & B[0];
  assign N[775] = A[8] & B[0];
  assign N[776] = N[663] & N[774];
  assign N[777] = N[666] & N[774];
  assign N[778] =  N[773] | N[776];
  assign N[779] = N[778] | N[777];
  assign N[780] = N[676] ^ N[673];
  assign N[781] = A[8] & B[1];
  assign N[782] = N[780] ^ N[781];
  assign N[783] = N[676] & N[673];
  assign N[784] = A[8] & B[1];
  assign N[785] = A[8] & B[1];
  assign N[786] = N[673] & N[784];
  assign N[787] = N[676] & N[784];
  assign N[788] =  N[783] | N[786];
  assign N[789] = N[788] | N[787];
  assign N[790] = N[686] ^ N[683];
  assign N[791] = A[8] & B[2];
  assign N[792] = N[790] ^ N[791];
  assign N[793] = N[686] & N[683];
  assign N[794] = A[8] & B[2];
  assign N[795] = A[8] & B[2];
  assign N[796] = N[683] & N[794];
  assign N[797] = N[686] & N[794];
  assign N[798] =  N[793] | N[796];
  assign N[799] = N[798] | N[797];
  assign N[800] = N[696] ^ N[693];
  assign N[801] = A[8] & B[3];
  assign N[802] = N[800] ^ N[801];
  assign N[803] = N[696] & N[693];
  assign N[804] = A[8] & B[3];
  assign N[805] = A[8] & B[3];
  assign N[806] = N[693] & N[804];
  assign N[807] = N[696] & N[804];
  assign N[808] =  N[803] | N[806];
  assign N[809] = N[808] | N[807];
  assign N[810] = N[706] ^ N[703];
  assign N[811] = A[8] & B[4];
  assign N[812] = N[810] ^ N[811];
  assign N[813] = N[706] & N[703];
  assign N[814] = A[8] & B[4];
  assign N[815] = A[8] & B[4];
  assign N[816] = N[703] & N[814];
  assign N[817] = N[706] & N[814];
  assign N[818] =  N[813] | N[816];
  assign N[819] = N[818] | N[817];
  assign N[820] = N[716] ^ N[713];
  assign N[821] = A[8] & B[5];
  assign N[822] = N[820] ^ N[821];
  assign N[823] = N[716] & N[713];
  assign N[824] = A[8] & B[5];
  assign N[825] = A[8] & B[5];
  assign N[826] = N[713] & N[824];
  assign N[827] = N[716] & N[824];
  assign N[828] =  N[823] | N[826];
  assign N[829] = N[828] | N[827];
  assign N[830] = N[726] ^ N[723];
  assign N[831] = A[8] & B[6];
  assign N[832] = N[830] ^ N[831];
  assign N[833] = N[726] & N[723];
  assign N[834] = A[8] & B[6];
  assign N[835] = A[8] & B[6];
  assign N[836] = N[723] & N[834];
  assign N[837] = N[726] & N[834];
  assign N[838] =  N[833] | N[836];
  assign N[839] = N[838] | N[837];
  assign N[840] = N[736] ^ N[733];
  assign N[841] = A[8] & B[7];
  assign N[842] = N[840] ^ N[841];
  assign N[843] = N[736] & N[733];
  assign N[844] = A[8] & B[7];
  assign N[845] = A[8] & B[7];
  assign N[846] = N[733] & N[844];
  assign N[847] = N[736] & N[844];
  assign N[848] =  N[843] | N[846];
  assign N[849] = N[848] | N[847];
  assign N[850] = N[746] ^ N[743];
  assign N[851] = A[8] & B[8];
  assign N[852] = N[850] ^ N[851];
  assign N[853] = N[746] & N[743];
  assign N[854] = A[8] & B[8];
  assign N[855] = A[8] & B[8];
  assign N[856] = N[743] & N[854];
  assign N[857] = N[746] & N[854];
  assign N[858] =  N[853] | N[856];
  assign N[859] = N[858] | N[857];
  assign N[860] = N[756] ^ N[753];
  assign N[861] = A[8] & B[9];
  assign N[862] = N[860] ^ N[861];
  assign N[863] = N[756] & N[753];
  assign N[864] = A[8] & B[9];
  assign N[865] = A[8] & B[9];
  assign N[866] = N[753] & N[864];
  assign N[867] = N[756] & N[864];
  assign N[868] =  N[863] | N[866];
  assign N[869] = N[868] | N[867];
  assign N[870] = N[766] ^ N[763];
  assign N[871] = A[8] & B[10];
  assign N[872] = N[870] ^ N[871];
  assign N[873] = N[766] & N[763];
  assign N[874] = A[8] & B[10];
  assign N[875] = A[8] & B[10];
  assign N[876] = N[763] & N[874];
  assign N[877] = N[766] & N[874];
  assign N[878] =  N[873] | N[876];
  assign N[879] = N[878] | N[877];
  assign N[880] = A[8] & B[11];
  assign N[881] = ~N[880];
  assign N[882] = N[769] ^  N[881];
  assign N[883] = A[8] & B[11];
  assign N[884] = ~N[883];
  assign N[885] = N[769] &  N[884];
  assign N[886] = N[782] ^ N[779];
  assign N[887] = A[9] & B[0];
  assign N[888] = N[886] ^ N[887];
  assign N[889] = N[782] & N[779];
  assign N[890] = A[9] & B[0];
  assign N[891] = A[9] & B[0];
  assign N[892] = N[779] & N[890];
  assign N[893] = N[782] & N[890];
  assign N[894] =  N[889] | N[892];
  assign N[895] = N[894] | N[893];
  assign N[896] = N[792] ^ N[789];
  assign N[897] = A[9] & B[1];
  assign N[898] = N[896] ^ N[897];
  assign N[899] = N[792] & N[789];
  assign N[900] = A[9] & B[1];
  assign N[901] = A[9] & B[1];
  assign N[902] = N[789] & N[900];
  assign N[903] = N[792] & N[900];
  assign N[904] =  N[899] | N[902];
  assign N[905] = N[904] | N[903];
  assign N[906] = N[802] ^ N[799];
  assign N[907] = A[9] & B[2];
  assign N[908] = N[906] ^ N[907];
  assign N[909] = N[802] & N[799];
  assign N[910] = A[9] & B[2];
  assign N[911] = A[9] & B[2];
  assign N[912] = N[799] & N[910];
  assign N[913] = N[802] & N[910];
  assign N[914] =  N[909] | N[912];
  assign N[915] = N[914] | N[913];
  assign N[916] = N[812] ^ N[809];
  assign N[917] = A[9] & B[3];
  assign N[918] = N[916] ^ N[917];
  assign N[919] = N[812] & N[809];
  assign N[920] = A[9] & B[3];
  assign N[921] = A[9] & B[3];
  assign N[922] = N[809] & N[920];
  assign N[923] = N[812] & N[920];
  assign N[924] =  N[919] | N[922];
  assign N[925] = N[924] | N[923];
  assign N[926] = N[822] ^ N[819];
  assign N[927] = A[9] & B[4];
  assign N[928] = N[926] ^ N[927];
  assign N[929] = N[822] & N[819];
  assign N[930] = A[9] & B[4];
  assign N[931] = A[9] & B[4];
  assign N[932] = N[819] & N[930];
  assign N[933] = N[822] & N[930];
  assign N[934] =  N[929] | N[932];
  assign N[935] = N[934] | N[933];
  assign N[936] = N[832] ^ N[829];
  assign N[937] = A[9] & B[5];
  assign N[938] = N[936] ^ N[937];
  assign N[939] = N[832] & N[829];
  assign N[940] = A[9] & B[5];
  assign N[941] = A[9] & B[5];
  assign N[942] = N[829] & N[940];
  assign N[943] = N[832] & N[940];
  assign N[944] =  N[939] | N[942];
  assign N[945] = N[944] | N[943];
  assign N[946] = N[842] ^ N[839];
  assign N[947] = A[9] & B[6];
  assign N[948] = N[946] ^ N[947];
  assign N[949] = N[842] & N[839];
  assign N[950] = A[9] & B[6];
  assign N[951] = A[9] & B[6];
  assign N[952] = N[839] & N[950];
  assign N[953] = N[842] & N[950];
  assign N[954] =  N[949] | N[952];
  assign N[955] = N[954] | N[953];
  assign N[956] = N[852] ^ N[849];
  assign N[957] = A[9] & B[7];
  assign N[958] = N[956] ^ N[957];
  assign N[959] = N[852] & N[849];
  assign N[960] = A[9] & B[7];
  assign N[961] = A[9] & B[7];
  assign N[962] = N[849] & N[960];
  assign N[963] = N[852] & N[960];
  assign N[964] =  N[959] | N[962];
  assign N[965] = N[964] | N[963];
  assign N[966] = N[862] ^ N[859];
  assign N[967] = A[9] & B[8];
  assign N[968] = N[966] ^ N[967];
  assign N[969] = N[862] & N[859];
  assign N[970] = A[9] & B[8];
  assign N[971] = A[9] & B[8];
  assign N[972] = N[859] & N[970];
  assign N[973] = N[862] & N[970];
  assign N[974] =  N[969] | N[972];
  assign N[975] = N[974] | N[973];
  assign N[976] = N[872] ^ N[869];
  assign N[977] = A[9] & B[9];
  assign N[978] = N[976] ^ N[977];
  assign N[979] = N[872] & N[869];
  assign N[980] = A[9] & B[9];
  assign N[981] = A[9] & B[9];
  assign N[982] = N[869] & N[980];
  assign N[983] = N[872] & N[980];
  assign N[984] =  N[979] | N[982];
  assign N[985] = N[984] | N[983];
  assign N[986] = N[882] ^ N[879];
  assign N[987] = A[9] & B[10];
  assign N[988] = N[986] ^ N[987];
  assign N[989] = N[882] & N[879];
  assign N[990] = A[9] & B[10];
  assign N[991] = A[9] & B[10];
  assign N[992] = N[879] & N[990];
  assign N[993] = N[882] & N[990];
  assign N[994] =  N[989] | N[992];
  assign N[995] = N[994] | N[993];
  assign N[996] = A[9] & B[11];
  assign N[997] = ~N[996];
  assign N[998] = N[885] ^  N[997];
  assign N[999] = A[9] & B[11];
  assign N[1000] = ~N[999];
  assign N[1001] = N[885] &  N[1000];
  assign N[1002] = N[898] ^ N[895];
  assign N[1003] = A[10] & B[0];
  assign N[1004] = N[1002] ^ N[1003];
  assign N[1005] = N[898] & N[895];
  assign N[1006] = A[10] & B[0];
  assign N[1007] = A[10] & B[0];
  assign N[1008] = N[895] & N[1006];
  assign N[1009] = N[898] & N[1006];
  assign N[1010] =  N[1005] | N[1008];
  assign N[1011] = N[1010] | N[1009];
  assign N[1012] = N[908] ^ N[905];
  assign N[1013] = A[10] & B[1];
  assign N[1014] = N[1012] ^ N[1013];
  assign N[1015] = N[908] & N[905];
  assign N[1016] = A[10] & B[1];
  assign N[1017] = A[10] & B[1];
  assign N[1018] = N[905] & N[1016];
  assign N[1019] = N[908] & N[1016];
  assign N[1020] =  N[1015] | N[1018];
  assign N[1021] = N[1020] | N[1019];
  assign N[1022] = N[918] ^ N[915];
  assign N[1023] = A[10] & B[2];
  assign N[1024] = N[1022] ^ N[1023];
  assign N[1025] = N[918] & N[915];
  assign N[1026] = A[10] & B[2];
  assign N[1027] = A[10] & B[2];
  assign N[1028] = N[915] & N[1026];
  assign N[1029] = N[918] & N[1026];
  assign N[1030] =  N[1025] | N[1028];
  assign N[1031] = N[1030] | N[1029];
  assign N[1032] = N[928] ^ N[925];
  assign N[1033] = A[10] & B[3];
  assign N[1034] = N[1032] ^ N[1033];
  assign N[1035] = N[928] & N[925];
  assign N[1036] = A[10] & B[3];
  assign N[1037] = A[10] & B[3];
  assign N[1038] = N[925] & N[1036];
  assign N[1039] = N[928] & N[1036];
  assign N[1040] =  N[1035] | N[1038];
  assign N[1041] = N[1040] | N[1039];
  assign N[1042] = N[938] ^ N[935];
  assign N[1043] = A[10] & B[4];
  assign N[1044] = N[1042] ^ N[1043];
  assign N[1045] = N[938] & N[935];
  assign N[1046] = A[10] & B[4];
  assign N[1047] = A[10] & B[4];
  assign N[1048] = N[935] & N[1046];
  assign N[1049] = N[938] & N[1046];
  assign N[1050] =  N[1045] | N[1048];
  assign N[1051] = N[1050] | N[1049];
  assign N[1052] = N[948] ^ N[945];
  assign N[1053] = A[10] & B[5];
  assign N[1054] = N[1052] ^ N[1053];
  assign N[1055] = N[948] & N[945];
  assign N[1056] = A[10] & B[5];
  assign N[1057] = A[10] & B[5];
  assign N[1058] = N[945] & N[1056];
  assign N[1059] = N[948] & N[1056];
  assign N[1060] =  N[1055] | N[1058];
  assign N[1061] = N[1060] | N[1059];
  assign N[1062] = N[958] ^ N[955];
  assign N[1063] = A[10] & B[6];
  assign N[1064] = N[1062] ^ N[1063];
  assign N[1065] = N[958] & N[955];
  assign N[1066] = A[10] & B[6];
  assign N[1067] = A[10] & B[6];
  assign N[1068] = N[955] & N[1066];
  assign N[1069] = N[958] & N[1066];
  assign N[1070] =  N[1065] | N[1068];
  assign N[1071] = N[1070] | N[1069];
  assign N[1072] = N[968] ^ N[965];
  assign N[1073] = A[10] & B[7];
  assign N[1074] = N[1072] ^ N[1073];
  assign N[1075] = N[968] & N[965];
  assign N[1076] = A[10] & B[7];
  assign N[1077] = A[10] & B[7];
  assign N[1078] = N[965] & N[1076];
  assign N[1079] = N[968] & N[1076];
  assign N[1080] =  N[1075] | N[1078];
  assign N[1081] = N[1080] | N[1079];
  assign N[1082] = N[978] ^ N[975];
  assign N[1083] = A[10] & B[8];
  assign N[1084] = N[1082] ^ N[1083];
  assign N[1085] = N[978] & N[975];
  assign N[1086] = A[10] & B[8];
  assign N[1087] = A[10] & B[8];
  assign N[1088] = N[975] & N[1086];
  assign N[1089] = N[978] & N[1086];
  assign N[1090] =  N[1085] | N[1088];
  assign N[1091] = N[1090] | N[1089];
  assign N[1092] = N[988] ^ N[985];
  assign N[1093] = A[10] & B[9];
  assign N[1094] = N[1092] ^ N[1093];
  assign N[1095] = N[988] & N[985];
  assign N[1096] = A[10] & B[9];
  assign N[1097] = A[10] & B[9];
  assign N[1098] = N[985] & N[1096];
  assign N[1099] = N[988] & N[1096];
  assign N[1100] =  N[1095] | N[1098];
  assign N[1101] = N[1100] | N[1099];
  assign N[1102] = N[998] ^ N[995];
  assign N[1103] = A[10] & B[10];
  assign N[1104] = N[1102] ^ N[1103];
  assign N[1105] = N[998] & N[995];
  assign N[1106] = A[10] & B[10];
  assign N[1107] = A[10] & B[10];
  assign N[1108] = N[995] & N[1106];
  assign N[1109] = N[998] & N[1106];
  assign N[1110] =  N[1105] | N[1108];
  assign N[1111] = N[1110] | N[1109];
  assign N[1112] = A[10] & B[11];
  assign N[1113] = ~N[1112];
  assign N[1114] = N[1001] ^  N[1113];
  assign N[1115] = A[10] & B[11];
  assign N[1116] = ~N[1115];
  assign N[1117] = N[1001] &  N[1116];
  assign N[1118] = N[1014] ^ N[1011];
  assign N[1119] = A[11] & B[0];
  assign N[1120] = ~N[1119];
  assign N[1121] = N[1118] ^  N[1120];
  assign N[1122] = N[1014] & N[1011];
  assign N[1123] = A[11] & B[0];
  assign N[1124] = A[11] & B[0];
  assign N[1125] = ~N[1123];
  assign N[1126] = N[1011] &  N[1125];
  assign N[1127] = ~N[1123];
  assign N[1128] = N[1014] &  N[1127];
  assign N[1129] =  N[1122] | N[1126];
  assign N[1130] = N[1129] | N[1128];
  assign N[1131] = N[1024] ^ N[1021];
  assign N[1132] = A[11] & B[1];
  assign N[1133] = ~N[1132];
  assign N[1134] = N[1131] ^  N[1133];
  assign N[1135] = N[1024] & N[1021];
  assign N[1136] = A[11] & B[1];
  assign N[1137] = A[11] & B[1];
  assign N[1138] = ~N[1136];
  assign N[1139] = N[1021] &  N[1138];
  assign N[1140] = ~N[1136];
  assign N[1141] = N[1024] &  N[1140];
  assign N[1142] =  N[1135] | N[1139];
  assign N[1143] = N[1142] | N[1141];
  assign N[1144] = N[1034] ^ N[1031];
  assign N[1145] = A[11] & B[2];
  assign N[1146] = ~N[1145];
  assign N[1147] = N[1144] ^  N[1146];
  assign N[1148] = N[1034] & N[1031];
  assign N[1149] = A[11] & B[2];
  assign N[1150] = A[11] & B[2];
  assign N[1151] = ~N[1149];
  assign N[1152] = N[1031] &  N[1151];
  assign N[1153] = ~N[1149];
  assign N[1154] = N[1034] &  N[1153];
  assign N[1155] =  N[1148] | N[1152];
  assign N[1156] = N[1155] | N[1154];
  assign N[1157] = N[1044] ^ N[1041];
  assign N[1158] = A[11] & B[3];
  assign N[1159] = ~N[1158];
  assign N[1160] = N[1157] ^  N[1159];
  assign N[1161] = N[1044] & N[1041];
  assign N[1162] = A[11] & B[3];
  assign N[1163] = A[11] & B[3];
  assign N[1164] = ~N[1162];
  assign N[1165] = N[1041] &  N[1164];
  assign N[1166] = ~N[1162];
  assign N[1167] = N[1044] &  N[1166];
  assign N[1168] =  N[1161] | N[1165];
  assign N[1169] = N[1168] | N[1167];
  assign N[1170] = N[1054] ^ N[1051];
  assign N[1171] = A[11] & B[4];
  assign N[1172] = ~N[1171];
  assign N[1173] = N[1170] ^  N[1172];
  assign N[1174] = N[1054] & N[1051];
  assign N[1175] = A[11] & B[4];
  assign N[1176] = A[11] & B[4];
  assign N[1177] = ~N[1175];
  assign N[1178] = N[1051] &  N[1177];
  assign N[1179] = ~N[1175];
  assign N[1180] = N[1054] &  N[1179];
  assign N[1181] =  N[1174] | N[1178];
  assign N[1182] = N[1181] | N[1180];
  assign N[1183] = N[1064] ^ N[1061];
  assign N[1184] = A[11] & B[5];
  assign N[1185] = ~N[1184];
  assign N[1186] = N[1183] ^  N[1185];
  assign N[1187] = N[1064] & N[1061];
  assign N[1188] = A[11] & B[5];
  assign N[1189] = A[11] & B[5];
  assign N[1190] = ~N[1188];
  assign N[1191] = N[1061] &  N[1190];
  assign N[1192] = ~N[1188];
  assign N[1193] = N[1064] &  N[1192];
  assign N[1194] =  N[1187] | N[1191];
  assign N[1195] = N[1194] | N[1193];
  assign N[1196] = N[1074] ^ N[1071];
  assign N[1197] = A[11] & B[6];
  assign N[1198] = ~N[1197];
  assign N[1199] = N[1196] ^  N[1198];
  assign N[1200] = N[1074] & N[1071];
  assign N[1201] = A[11] & B[6];
  assign N[1202] = A[11] & B[6];
  assign N[1203] = ~N[1201];
  assign N[1204] = N[1071] &  N[1203];
  assign N[1205] = ~N[1201];
  assign N[1206] = N[1074] &  N[1205];
  assign N[1207] =  N[1200] | N[1204];
  assign N[1208] = N[1207] | N[1206];
  assign N[1209] = N[1084] ^ N[1081];
  assign N[1210] = A[11] & B[7];
  assign N[1211] = ~N[1210];
  assign N[1212] = N[1209] ^  N[1211];
  assign N[1213] = N[1084] & N[1081];
  assign N[1214] = A[11] & B[7];
  assign N[1215] = A[11] & B[7];
  assign N[1216] = ~N[1214];
  assign N[1217] = N[1081] &  N[1216];
  assign N[1218] = ~N[1214];
  assign N[1219] = N[1084] &  N[1218];
  assign N[1220] =  N[1213] | N[1217];
  assign N[1221] = N[1220] | N[1219];
  assign N[1222] = N[1094] ^ N[1091];
  assign N[1223] = A[11] & B[8];
  assign N[1224] = ~N[1223];
  assign N[1225] = N[1222] ^  N[1224];
  assign N[1226] = N[1094] & N[1091];
  assign N[1227] = A[11] & B[8];
  assign N[1228] = A[11] & B[8];
  assign N[1229] = ~N[1227];
  assign N[1230] = N[1091] &  N[1229];
  assign N[1231] = ~N[1227];
  assign N[1232] = N[1094] &  N[1231];
  assign N[1233] =  N[1226] | N[1230];
  assign N[1234] = N[1233] | N[1232];
  assign N[1235] = N[1104] ^ N[1101];
  assign N[1236] = A[11] & B[9];
  assign N[1237] = ~N[1236];
  assign N[1238] = N[1235] ^  N[1237];
  assign N[1239] = N[1104] & N[1101];
  assign N[1240] = A[11] & B[9];
  assign N[1241] = A[11] & B[9];
  assign N[1242] = ~N[1240];
  assign N[1243] = N[1101] &  N[1242];
  assign N[1244] = ~N[1240];
  assign N[1245] = N[1104] &  N[1244];
  assign N[1246] =  N[1239] | N[1243];
  assign N[1247] = N[1246] | N[1245];
  assign N[1248] = N[1114] ^ N[1111];
  assign N[1249] = A[11] & B[10];
  assign N[1250] = ~N[1249];
  assign N[1251] = N[1248] ^  N[1250];
  assign N[1252] = N[1114] & N[1111];
  assign N[1253] = A[11] & B[10];
  assign N[1254] = A[11] & B[10];
  assign N[1255] = ~N[1253];
  assign N[1256] = N[1111] &  N[1255];
  assign N[1257] = ~N[1253];
  assign N[1258] = N[1114] &  N[1257];
  assign N[1259] =  N[1252] | N[1256];
  assign N[1260] = N[1259] | N[1258];
  assign N[1261] = A[11] & B[11];
  assign N[1262] = N[1117] ^ N[1261];
  assign N[1263] = A[11] & B[11];
  assign N[1264] = N[1117] & N[1263];
  assign N[1265] = N[1134] ^ N[1130];
  assign N[1266] = N[1134] & N[1130];
  assign N[1267] = N[1147] ^ N[1266];
  assign N[1268] = N[1267] ^ N[1143];
  assign N[1269] = N[1147] & N[1266];
  assign N[1270] = N[1266] & N[1143];
  assign N[1271] = N[1147] & N[1143];
  assign N[1272] =  N[1269] | N[1270];
  assign N[1273] = N[1272] | N[1271];
  assign N[1274] = N[1160] ^ N[1273];
  assign N[1275] = N[1274] ^ N[1156];
  assign N[1276] = N[1160] & N[1273];
  assign N[1277] = N[1273] & N[1156];
  assign N[1278] = N[1160] & N[1156];
  assign N[1279] =  N[1276] | N[1277];
  assign N[1280] = N[1279] | N[1278];
  assign N[1281] = N[1173] ^ N[1280];
  assign N[1282] = N[1281] ^ N[1169];
  assign N[1283] = N[1173] & N[1280];
  assign N[1284] = N[1280] & N[1169];
  assign N[1285] = N[1173] & N[1169];
  assign N[1286] =  N[1283] | N[1284];
  assign N[1287] = N[1286] | N[1285];
  assign N[1288] = N[1186] ^ N[1287];
  assign N[1289] = N[1288] ^ N[1182];
  assign N[1290] = N[1186] & N[1287];
  assign N[1291] = N[1287] & N[1182];
  assign N[1292] = N[1186] & N[1182];
  assign N[1293] =  N[1290] | N[1291];
  assign N[1294] = N[1293] | N[1292];
  assign N[1295] = N[1199] ^ N[1294];
  assign N[1296] = N[1295] ^ N[1195];
  assign N[1297] = N[1199] & N[1294];
  assign N[1298] = N[1294] & N[1195];
  assign N[1299] = N[1199] & N[1195];
  assign N[1300] =  N[1297] | N[1298];
  assign N[1301] = N[1300] | N[1299];
  assign N[1302] = N[1212] ^ N[1301];
  assign N[1303] = N[1302] ^ N[1208];
  assign N[1304] = N[1212] & N[1301];
  assign N[1305] = N[1301] & N[1208];
  assign N[1306] = N[1212] & N[1208];
  assign N[1307] =  N[1304] | N[1305];
  assign N[1308] = N[1307] | N[1306];
  assign N[1309] = N[1225] ^ N[1308];
  assign N[1310] = N[1309] ^ N[1221];
  assign N[1311] = N[1225] & N[1308];
  assign N[1312] = N[1308] & N[1221];
  assign N[1313] = N[1225] & N[1221];
  assign N[1314] =  N[1311] | N[1312];
  assign N[1315] = N[1314] | N[1313];
  assign N[1316] = N[1238] ^ N[1315];
  assign N[1317] = N[1316] ^ N[1234];
  assign N[1318] = N[1238] & N[1315];
  assign N[1319] = N[1315] & N[1234];
  assign N[1320] = N[1238] & N[1234];
  assign N[1321] =  N[1318] | N[1319];
  assign N[1322] = N[1321] | N[1320];
  assign N[1323] = N[1251] ^ N[1322];
  assign N[1324] = N[1323] ^ N[1247];
  assign N[1325] = N[1251] & N[1322];
  assign N[1326] = N[1322] & N[1247];
  assign N[1327] = N[1251] & N[1247];
  assign N[1328] =  N[1325] | N[1326];
  assign N[1329] = N[1328] | N[1327];
  assign N[1330] = N[1262] ^ N[1329];
  assign N[1331] = N[1330] ^ N[1260];
  assign N[1332] = N[1262] & N[1329];
  assign N[1333] = N[1329] & N[1260];
  assign N[1334] = N[1262] & N[1260];
  assign N[1335] =  N[1332] | N[1333];
  assign N[1336] = N[1335] | N[1334];
  assign N[1337] = 1'b1 ^ N[1336];
  assign N[1338] = N[1337] ^ N[1264];
  assign N[1339] = 1'b1 & N[1336];
  assign N[1340] = N[1336] & N[1264];
  assign N[1341] = 1'b1 & N[1264];
  assign N[1342] =  N[1339] | N[1340];
  assign N[1343] = N[1342] | N[1341];
  assign O = {N[1338],N[1331],N[1324],N[1317],N[1310],N[1303],N[1296],N[1289],N[1282],N[1275],N[1268],N[1265],N[1121],N[1004],N[888],N[772],N[656],N[540],N[424],N[308],N[192],N[76],N[25],N[1]};

endmodule